*mosfet
.model nmos_intr nmos level=1 kp=50u vto=0.5 lambda=0.1 gamma=0.6 phi=0.8 tox=150n cgdo=0 cgso=0
vgs  1  0 dc 1.25
vds  2 0  dc 1

*   drain gate source bulk
mn1  2 1 0 0 nmos_intr w=.2u 
.dc vgs 1 3.3 0.5 vds 1 3.3 0.5 

.control
     run 
      save @mn1[w]
     
      print v(2) i(vds) @mn1[w]


      
     



  
    
.endc

.end
